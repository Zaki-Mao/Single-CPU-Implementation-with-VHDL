----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:23:48 05/18/2021 
-- Design Name: 
-- Module Name:    jumpaddressshift - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity myjas16 is
port(
	input : in STD_LOGIC_VECTOR(27 downto 0);
	output : out STD_LOGIC_VECTOR(27 downto 0)); 
end myjas16;

architecture Behavioral of myjas16 is

begin
	output <= to_STDLOGICVECTOR(to_bitvector(input) sla 2);

end Behavioral;
